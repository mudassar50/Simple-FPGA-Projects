module ALU2Bit( // @[:@3.2]
  input        clock, // @[:@4.4]
  input        reset, // @[:@5.4]
  input  [1:0] io_A, // @[:@6.4]
  input  [1:0] io_B, // @[:@6.4]
  input  [1:0] io_Op, // @[:@6.4]
  output [1:0] io_Result, // @[:@6.4]
  output [3:0] io_LED // @[:@6.4]
);
  wire [2:0] _T_17; // @[2bitAlu.scala 17:23:@8.4]
  wire [1:0] _T_18; // @[2bitAlu.scala 17:23:@9.4]
  wire [2:0] _T_20; // @[2bitAlu.scala 18:23:@10.4]
  wire [2:0] _T_21; // @[2bitAlu.scala 18:23:@11.4]
  wire [1:0] _T_22; // @[2bitAlu.scala 18:23:@12.4]
  wire [1:0] _T_24; // @[2bitAlu.scala 19:23:@13.4]
  wire [1:0] _T_26; // @[2bitAlu.scala 20:23:@14.4]
  wire  _T_27; // @[Mux.scala 46:19:@15.4]
  wire [1:0] _T_28; // @[Mux.scala 46:16:@16.4]
  wire  _T_29; // @[Mux.scala 46:19:@17.4]
  wire [1:0] _T_30; // @[Mux.scala 46:16:@18.4]
  wire  _T_31; // @[Mux.scala 46:19:@19.4]
  wire [1:0] _T_32; // @[Mux.scala 46:16:@20.4]
  wire  _T_33; // @[Mux.scala 46:19:@21.4]
  assign _T_17 = io_A + io_B; // @[2bitAlu.scala 17:23:@8.4]
  assign _T_18 = io_A + io_B; // @[2bitAlu.scala 17:23:@9.4]
  assign _T_20 = io_A - io_B; // @[2bitAlu.scala 18:23:@10.4]
  assign _T_21 = $unsigned(_T_20); // @[2bitAlu.scala 18:23:@11.4]
  assign _T_22 = _T_21[1:0]; // @[2bitAlu.scala 18:23:@12.4]
  assign _T_24 = io_A & io_B; // @[2bitAlu.scala 19:23:@13.4]
  assign _T_26 = io_A | io_B; // @[2bitAlu.scala 20:23:@14.4]
  assign _T_27 = 2'h3 == io_Op; // @[Mux.scala 46:19:@15.4]
  assign _T_28 = _T_27 ? _T_26 : 2'h0; // @[Mux.scala 46:16:@16.4]
  assign _T_29 = 2'h2 == io_Op; // @[Mux.scala 46:19:@17.4]
  assign _T_30 = _T_29 ? _T_24 : _T_28; // @[Mux.scala 46:16:@18.4]
  assign _T_31 = 2'h1 == io_Op; // @[Mux.scala 46:19:@19.4]
  assign _T_32 = _T_31 ? _T_22 : _T_30; // @[Mux.scala 46:16:@20.4]
  assign _T_33 = 2'h0 == io_Op; // @[Mux.scala 46:19:@21.4]
  assign io_Result = _T_33 ? _T_18 : _T_32; // @[2bitAlu.scala 16:13:@23.4]
  assign io_LED = {2'h0,io_Result}; // @[2bitAlu.scala 24:10:@25.4]
endmodule
